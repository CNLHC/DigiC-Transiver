// OFDM_Modulation.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module OFDM_Modulation (
		input  wire        clk_clk,                     //           clk.clk
		input  wire        fft_ii_0_sink_valid,         // fft_ii_0_sink.valid
		output wire        fft_ii_0_sink_ready,         //              .ready
		input  wire [1:0]  fft_ii_0_sink_error,         //              .error
		input  wire        fft_ii_0_sink_startofpacket, //              .startofpacket
		input  wire        fft_ii_0_sink_endofpacket,   //              .endofpacket
		input  wire [32:0] fft_ii_0_sink_data,          //              .data
		input  wire        reset_reset_n                //         reset.reset_n
	);

	wire         fft_ii_0_source_valid;                 // fft_ii_0:source_valid -> avalon_st_adapter:in_0_valid
	wire  [37:0] fft_ii_0_source_data;                  // fft_ii_0:source_data -> avalon_st_adapter:in_0_data
	wire         fft_ii_0_source_ready;                 // avalon_st_adapter:in_0_ready -> fft_ii_0:source_ready
	wire         fft_ii_0_source_startofpacket;         // fft_ii_0:source_sop -> avalon_st_adapter:in_0_startofpacket
	wire   [1:0] fft_ii_0_source_error;                 // fft_ii_0:source_error -> avalon_st_adapter:in_0_error
	wire         fft_ii_0_source_endofpacket;           // fft_ii_0:source_eop -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;         // avalon_st_adapter:out_0_valid -> OFDM_Cyclic_Prefix_Adder_0:asi_in0_valid
	wire  [37:0] avalon_st_adapter_out_0_data;          // avalon_st_adapter:out_0_data -> OFDM_Cyclic_Prefix_Adder_0:asi_in0_data
	wire         avalon_st_adapter_out_0_ready;         // OFDM_Cyclic_Prefix_Adder_0:asi_in0_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket; // avalon_st_adapter:out_0_startofpacket -> OFDM_Cyclic_Prefix_Adder_0:asi_in0_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;   // avalon_st_adapter:out_0_endofpacket -> OFDM_Cyclic_Prefix_Adder_0:asi_in0_endofpacket
	wire         rst_controller_reset_out_reset;        // rst_controller:reset_out -> [OFDM_Cyclic_Prefix_Adder_0:reset_reset, avalon_st_adapter:in_rst_0_reset, fft_ii_0:reset_n]
	wire  [15:0] fft_ii_0_source_imag;                  // port fragment
	wire  [15:0] fft_ii_0_source_real;                  // port fragment
	wire   [5:0] fft_ii_0_source_exp;                   // port fragment

	OFDM_Cyclic_Prefix_Adder #(
		.Packet_Length (1024),
		.CP_Length     (128)
	) ofdm_cyclic_prefix_adder_0 (
		.asi_in0_data           (avalon_st_adapter_out_0_data),          //  asi_in0.data
		.asi_in0_ready          (avalon_st_adapter_out_0_ready),         //         .ready
		.asi_in0_valid          (avalon_st_adapter_out_0_valid),         //         .valid
		.asi_in0_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.asi_in0_startofpacket  (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.clock_clk              (clk_clk),                               //    clock.clk
		.reset_reset            (rst_controller_reset_out_reset),        //    reset.reset
		.aso_out0_data          (),                                      // aso_out0.data
		.aso_out0_ready         (),                                      //         .ready
		.aso_out0_valid         (),                                      //         .valid
		.aso_out0_endofpacket   (),                                      //         .endofpacket
		.aso_out0_startofpacket ()                                       //         .startofpacket
	);

	OFDM_Modulation_fft_ii_0 fft_ii_0 (
		.clk          (clk_clk),                         //    clk.clk
		.reset_n      (~rst_controller_reset_out_reset), //    rst.reset_n
		.sink_valid   (fft_ii_0_sink_valid),             //   sink.valid
		.sink_ready   (fft_ii_0_sink_ready),             //       .ready
		.sink_error   (fft_ii_0_sink_error),             //       .error
		.sink_sop     (fft_ii_0_sink_startofpacket),     //       .startofpacket
		.sink_eop     (fft_ii_0_sink_endofpacket),       //       .endofpacket
		.sink_real    (fft_ii_0_sink_data[32:17]),       //       .data
		.sink_imag    (fft_ii_0_sink_data[16:1]),        //       .data
		.inverse      (fft_ii_0_sink_data[0]),           //       .data
		.source_valid (fft_ii_0_source_valid),           // source.valid
		.source_ready (fft_ii_0_source_ready),           //       .ready
		.source_error (fft_ii_0_source_error),           //       .error
		.source_sop   (fft_ii_0_source_startofpacket),   //       .startofpacket
		.source_eop   (fft_ii_0_source_endofpacket),     //       .endofpacket
		.source_real  (fft_ii_0_source_real[15:0]),      //       .data
		.source_imag  (fft_ii_0_source_imag[15:0]),      //       .data
		.source_exp   (fft_ii_0_source_exp[5:0])         //       .data
	);

	OFDM_Modulation_avalon_st_adapter #(
		.inBitsPerSymbol (38),
		.inUsePackets    (1),
		.inDataWidth     (38),
		.inChannelWidth  (0),
		.inErrorWidth    (2),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (38),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (fft_ii_0_source_data),                  //     in_0.data
		.in_0_valid          (fft_ii_0_source_valid),                 //         .valid
		.in_0_ready          (fft_ii_0_source_ready),                 //         .ready
		.in_0_startofpacket  (fft_ii_0_source_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (fft_ii_0_source_endofpacket),           //         .endofpacket
		.in_0_error          (fft_ii_0_source_error),                 //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)    //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	assign fft_ii_0_source_data = { fft_ii_0_source_real[15:0], fft_ii_0_source_imag[15:0], fft_ii_0_source_exp[5:0] };

endmodule
