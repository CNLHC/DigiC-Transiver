// DigiCQSysTop_DigiCQSys_0.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module DigiCQSysTop_DigiCQSys_0 (
		input  wire        global_reset_reset_n,                    //              global_reset.reset_n
		output wire        pll_0_locked_export,                     //              pll_0_locked.export
		output wire        pll_0_outclk_1_clk,                      //            pll_0_outclk_1.clk
		output wire        pll_0_outclk_10_clk,                     //           pll_0_outclk_10.clk
		output wire        pll_0_outclk_120_clk,                    //          pll_0_outclk_120.clk
		output wire        pll_0_outclk_20_clk,                     //           pll_0_outclk_20.clk
		input  wire        pll_0_refclk_clk,                        //              pll_0_refclk.clk
		output wire [32:0] qam_modulation_0_aso_out0_data,          // qam_modulation_0_aso_out0.data
		input  wire        qam_modulation_0_aso_out0_ready,         //                          .ready
		output wire        qam_modulation_0_aso_out0_valid,         //                          .valid
		output wire        qam_modulation_0_aso_out0_empty,         //                          .empty
		output wire        qam_modulation_0_aso_out0_endofpacket,   //                          .endofpacket
		output wire        qam_modulation_0_aso_out0_startofpacket, //                          .startofpacket
		input  wire        qsys_clkin_clk,                          //                qsys_clkin.clk
		input  wire        spislave_0_export_0_mosi,                //       spislave_0_export_0.mosi
		input  wire        spislave_0_export_0_nss,                 //                          .nss
		inout  wire        spislave_0_export_0_miso,                //                          .miso
		input  wire        spislave_0_export_0_sclk                 //                          .sclk
	);

	wire         spislave_0_avalon_streaming_source_valid;               // spislave_0:stsourcevalid -> st_bytes_to_packets_0:in_valid
	wire   [7:0] spislave_0_avalon_streaming_source_data;                // spislave_0:stsourcedata -> st_bytes_to_packets_0:in_data
	wire         spislave_0_avalon_streaming_source_ready;               // st_bytes_to_packets_0:in_ready -> spislave_0:stsourceready
	wire         st_bytes_to_packets_0_out_packets_stream_valid;         // st_bytes_to_packets_0:out_valid -> avalon_st_adapter:in_0_valid
	wire   [7:0] st_bytes_to_packets_0_out_packets_stream_data;          // st_bytes_to_packets_0:out_data -> avalon_st_adapter:in_0_data
	wire         st_bytes_to_packets_0_out_packets_stream_ready;         // avalon_st_adapter:in_0_ready -> st_bytes_to_packets_0:out_ready
	wire   [7:0] st_bytes_to_packets_0_out_packets_stream_channel;       // st_bytes_to_packets_0:out_channel -> avalon_st_adapter:in_0_channel
	wire         st_bytes_to_packets_0_out_packets_stream_startofpacket; // st_bytes_to_packets_0:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         st_bytes_to_packets_0_out_packets_stream_endofpacket;   // st_bytes_to_packets_0:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                          // avalon_st_adapter:out_0_valid -> QAM_Modulation_0:asi_in0_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                           // avalon_st_adapter:out_0_data -> QAM_Modulation_0:asi_in0_data
	wire         avalon_st_adapter_out_0_ready;                          // QAM_Modulation_0:asi_in0_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                  // avalon_st_adapter:out_0_startofpacket -> QAM_Modulation_0:asi_in0_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                    // avalon_st_adapter:out_0_endofpacket -> QAM_Modulation_0:asi_in0_endofpacket
	wire   [1:0] avalon_st_adapter_out_0_empty;                          // avalon_st_adapter:out_0_empty -> QAM_Modulation_0:asi_in0_empty
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [QAM_Modulation_0:reset_reset, avalon_st_adapter:in_rst_0_reset, spislave_0:nreset, st_bytes_to_packets_0:reset_n]

	QAM_Modulation #(
		.PACKET_LENGTH (1024)
	) qam_modulation_0 (
		.asi_in0_data           (avalon_st_adapter_out_0_data),            //  asi_in0.data
		.asi_in0_ready          (avalon_st_adapter_out_0_ready),           //         .ready
		.asi_in0_valid          (avalon_st_adapter_out_0_valid),           //         .valid
		.asi_in0_startofpacket  (avalon_st_adapter_out_0_startofpacket),   //         .startofpacket
		.asi_in0_endofpacket    (avalon_st_adapter_out_0_endofpacket),     //         .endofpacket
		.asi_in0_empty          (avalon_st_adapter_out_0_empty),           //         .empty
		.clock_clk              (qsys_clkin_clk),                          //    clock.clk
		.reset_reset            (rst_controller_reset_out_reset),          //    reset.reset
		.aso_out0_data          (qam_modulation_0_aso_out0_data),          // aso_out0.data
		.aso_out0_ready         (qam_modulation_0_aso_out0_ready),         //         .ready
		.aso_out0_valid         (qam_modulation_0_aso_out0_valid),         //         .valid
		.aso_out0_empty         (qam_modulation_0_aso_out0_empty),         //         .empty
		.aso_out0_endofpacket   (qam_modulation_0_aso_out0_endofpacket),   //         .endofpacket
		.aso_out0_startofpacket (qam_modulation_0_aso_out0_startofpacket)  //         .startofpacket
	);

	DigiCQSysTop_DigiCQSys_0_pll_0 pll_0 (
		.refclk   (pll_0_refclk_clk),      //  refclk.clk
		.rst      (~global_reset_reset_n), //   reset.reset
		.outclk_0 (pll_0_outclk_1_clk),    // outclk0.clk
		.outclk_1 (pll_0_outclk_10_clk),   // outclk1.clk
		.outclk_2 (pll_0_outclk_20_clk),   // outclk2.clk
		.outclk_3 (pll_0_outclk_120_clk),  // outclk3.clk
		.locked   (pll_0_locked_export)    //  locked.export
	);

	SPIPhy #(
		.SYNC_DEPTH (2)
	) spislave_0 (
		.sysclk        (qsys_clkin_clk),                           //              clock_sink.clk
		.nreset        (~rst_controller_reset_out_reset),          //        clock_sink_reset.reset_n
		.mosi          (spislave_0_export_0_mosi),                 //                export_0.export
		.nss           (spislave_0_export_0_nss),                  //                        .export
		.miso          (spislave_0_export_0_miso),                 //                        .export
		.sclk          (spislave_0_export_0_sclk),                 //                        .export
		.stsourceready (spislave_0_avalon_streaming_source_ready), // avalon_streaming_source.ready
		.stsourcevalid (spislave_0_avalon_streaming_source_valid), //                        .valid
		.stsourcedata  (spislave_0_avalon_streaming_source_data),  //                        .data
		.stsinkvalid   (),                                         //   avalon_streaming_sink.valid
		.stsinkdata    (),                                         //                        .data
		.stsinkready   ()                                          //                        .ready
	);

	altera_avalon_st_bytes_to_packets #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) st_bytes_to_packets_0 (
		.clk               (qsys_clkin_clk),                                         //                clk.clk
		.reset_n           (~rst_controller_reset_out_reset),                        //          clk_reset.reset_n
		.out_channel       (st_bytes_to_packets_0_out_packets_stream_channel),       // out_packets_stream.channel
		.out_ready         (st_bytes_to_packets_0_out_packets_stream_ready),         //                   .ready
		.out_valid         (st_bytes_to_packets_0_out_packets_stream_valid),         //                   .valid
		.out_data          (st_bytes_to_packets_0_out_packets_stream_data),          //                   .data
		.out_startofpacket (st_bytes_to_packets_0_out_packets_stream_startofpacket), //                   .startofpacket
		.out_endofpacket   (st_bytes_to_packets_0_out_packets_stream_endofpacket),   //                   .endofpacket
		.in_ready          (spislave_0_avalon_streaming_source_ready),               //    in_bytes_stream.ready
		.in_valid          (spislave_0_avalon_streaming_source_valid),               //                   .valid
		.in_data           (spislave_0_avalon_streaming_source_data)                 //                   .data
	);

	DigiCQSysTop_DigiCQSys_0_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (8),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (qsys_clkin_clk),                                         // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                         // in_rst_0.reset
		.in_0_data           (st_bytes_to_packets_0_out_packets_stream_data),          //     in_0.data
		.in_0_valid          (st_bytes_to_packets_0_out_packets_stream_valid),         //         .valid
		.in_0_ready          (st_bytes_to_packets_0_out_packets_stream_ready),         //         .ready
		.in_0_startofpacket  (st_bytes_to_packets_0_out_packets_stream_startofpacket), //         .startofpacket
		.in_0_endofpacket    (st_bytes_to_packets_0_out_packets_stream_endofpacket),   //         .endofpacket
		.in_0_channel        (st_bytes_to_packets_0_out_packets_stream_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                           //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                          //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                          //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),                    //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)                           //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~global_reset_reset_n),          // reset_in0.reset
		.clk            (qsys_clkin_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
