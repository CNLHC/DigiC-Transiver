
module DigiCQSys (
	global_reset_reset_n,
	qsys_clkin_clk,
	receivertopqsys_0_ofdmadccontrol_external_adc_RealData,
	receivertopqsys_0_ofdmadccontrol_external_adc_ImagData,
	signaltaopll_outclk0_clk,
	systemclockpll_addaclk_clk,
	transmittertopqsys_0_externalspi_export_0_mosi,
	transmittertopqsys_0_externalspi_export_0_nss,
	transmittertopqsys_0_externalspi_export_0_miso,
	transmittertopqsys_0_externalspi_export_0_sclk,
	transmittertopqsys_0_ofdmdaccontrol_dac_control_chadata,
	transmittertopqsys_0_ofdmdaccontrol_dac_control_chbdata);	

	input		global_reset_reset_n;
	input		qsys_clkin_clk;
	input	[13:0]	receivertopqsys_0_ofdmadccontrol_external_adc_RealData;
	input	[13:0]	receivertopqsys_0_ofdmadccontrol_external_adc_ImagData;
	output		signaltaopll_outclk0_clk;
	output		systemclockpll_addaclk_clk;
	input		transmittertopqsys_0_externalspi_export_0_mosi;
	input		transmittertopqsys_0_externalspi_export_0_nss;
	inout		transmittertopqsys_0_externalspi_export_0_miso;
	input		transmittertopqsys_0_externalspi_export_0_sclk;
	output	[13:0]	transmittertopqsys_0_ofdmdaccontrol_dac_control_chadata;
	output	[13:0]	transmittertopqsys_0_ofdmdaccontrol_dac_control_chbdata;
endmodule
