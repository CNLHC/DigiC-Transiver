// OFDMCPAdder.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module OFDMCPAdder (
		input  wire [21:0] avalon_st_demux_0_asi_in0_data,          // avalon_st_demux_0_asi_in0.data
		output wire        avalon_st_demux_0_asi_in0_ready,         //                          .ready
		input  wire        avalon_st_demux_0_asi_in0_valid,         //                          .valid
		input  wire        avalon_st_demux_0_asi_in0_endofpacket,   //                          .endofpacket
		input  wire        avalon_st_demux_0_asi_in0_startofpacket, //                          .startofpacket
		input  wire        clk_clk,                                 //                       clk.clk
		output wire [21:0] cpadderrouter_0_data_out_data,           //  cpadderrouter_0_data_out.data
		output wire        cpadderrouter_0_data_out_valid,          //                          .valid
		output wire [1:0]  cpadderrouter_0_data_out_error,          //                          .error
		output wire        cpadderrouter_0_data_out_endofpacket,    //                          .endofpacket
		output wire        cpadderrouter_0_data_out_startofpacket,  //                          .startofpacket
		input  wire        reset_reset_n                            //                     reset.reset_n
	);

	wire         avalon_st_demux_0_aso_out0_valid;         // Avalon_ST_Demux_0:aso_out0_valid -> CPAdderRouter_0:asi_in0_valid
	wire  [21:0] avalon_st_demux_0_aso_out0_data;          // Avalon_ST_Demux_0:aso_out0_data -> CPAdderRouter_0:asi_in0_data
	wire         avalon_st_demux_0_aso_out0_ready;         // CPAdderRouter_0:asi_in0_ready -> Avalon_ST_Demux_0:aso_out0_ready
	wire         avalon_st_demux_0_aso_out0_startofpacket; // Avalon_ST_Demux_0:aso_out0_startofpacket -> CPAdderRouter_0:asi_in0_startofpacket
	wire         avalon_st_demux_0_aso_out0_endofpacket;   // Avalon_ST_Demux_0:aso_out0_endofpacket -> CPAdderRouter_0:asi_in0_endofpacket
	wire         avalon_st_demux_0_aso_out1_valid;         // Avalon_ST_Demux_0:aso_out1_valid -> sc_fifo_0:in_valid
	wire  [21:0] avalon_st_demux_0_aso_out1_data;          // Avalon_ST_Demux_0:aso_out1_data -> sc_fifo_0:in_data
	wire         avalon_st_demux_0_aso_out1_ready;         // sc_fifo_0:in_ready -> Avalon_ST_Demux_0:aso_out1_ready
	wire         avalon_st_demux_0_aso_out1_startofpacket; // Avalon_ST_Demux_0:aso_out1_startofpacket -> sc_fifo_0:in_startofpacket
	wire         avalon_st_demux_0_aso_out1_endofpacket;   // Avalon_ST_Demux_0:aso_out1_endofpacket -> sc_fifo_0:in_endofpacket
	wire         sc_fifo_0_out_valid;                      // sc_fifo_0:out_valid -> CPAdderRouter_0:buffer_in_valid
	wire  [21:0] sc_fifo_0_out_data;                       // sc_fifo_0:out_data -> CPAdderRouter_0:buffer_in_data
	wire         sc_fifo_0_out_ready;                      // CPAdderRouter_0:buffer_in_ready -> sc_fifo_0:out_ready
	wire         sc_fifo_0_out_startofpacket;              // sc_fifo_0:out_startofpacket -> CPAdderRouter_0:buffer_in_startofpacket
	wire         sc_fifo_0_out_endofpacket;                // sc_fifo_0:out_endofpacket -> CPAdderRouter_0:buffer_in_endofpacket
	wire         rst_controller_reset_out_reset;           // rst_controller:reset_out -> [Avalon_ST_Demux_0:reset_reset, CPAdderRouter_0:reset_reset, sc_fifo_0:reset]

	Avalon_ST_Demux avalon_st_demux_0 (
		.asi_in0_data           (avalon_st_demux_0_asi_in0_data),           //  asi_in0.data
		.asi_in0_ready          (avalon_st_demux_0_asi_in0_ready),          //         .ready
		.asi_in0_valid          (avalon_st_demux_0_asi_in0_valid),          //         .valid
		.asi_in0_endofpacket    (avalon_st_demux_0_asi_in0_endofpacket),    //         .endofpacket
		.asi_in0_startofpacket  (avalon_st_demux_0_asi_in0_startofpacket),  //         .startofpacket
		.clock_clk              (clk_clk),                                  //    clock.clk
		.reset_reset            (rst_controller_reset_out_reset),           //    reset.reset
		.aso_out0_data          (avalon_st_demux_0_aso_out0_data),          // aso_out0.data
		.aso_out0_ready         (avalon_st_demux_0_aso_out0_ready),         //         .ready
		.aso_out0_valid         (avalon_st_demux_0_aso_out0_valid),         //         .valid
		.aso_out0_endofpacket   (avalon_st_demux_0_aso_out0_endofpacket),   //         .endofpacket
		.aso_out0_startofpacket (avalon_st_demux_0_aso_out0_startofpacket), //         .startofpacket
		.aso_out1_data          (avalon_st_demux_0_aso_out1_data),          // aso_out1.data
		.aso_out1_ready         (avalon_st_demux_0_aso_out1_ready),         //         .ready
		.aso_out1_valid         (avalon_st_demux_0_aso_out1_valid),         //         .valid
		.aso_out1_endofpacket   (avalon_st_demux_0_aso_out1_endofpacket),   //         .endofpacket
		.aso_out1_startofpacket (avalon_st_demux_0_aso_out1_startofpacket)  //         .startofpacket
	);

	OFDM_Cyclic_Prefix_Adder #(
		.Packet_Length (1024),
		.CP_Length     (256)
	) cpadderrouter_0 (
		.asi_in0_data            (avalon_st_demux_0_aso_out0_data),          //   asi_in0.data
		.asi_in0_valid           (avalon_st_demux_0_aso_out0_valid),         //          .valid
		.asi_in0_endofpacket     (avalon_st_demux_0_aso_out0_endofpacket),   //          .endofpacket
		.asi_in0_startofpacket   (avalon_st_demux_0_aso_out0_startofpacket), //          .startofpacket
		.asi_in0_ready           (avalon_st_demux_0_aso_out0_ready),         //          .ready
		.clock_clk               (clk_clk),                                  //     clock.clk
		.reset_reset             (rst_controller_reset_out_reset),           //     reset.reset
		.buffer_in_data          (sc_fifo_0_out_data),                       // buffer_in.data
		.buffer_in_ready         (sc_fifo_0_out_ready),                      //          .ready
		.buffer_in_valid         (sc_fifo_0_out_valid),                      //          .valid
		.buffer_in_startofpacket (sc_fifo_0_out_startofpacket),              //          .startofpacket
		.buffer_in_endofpacket   (sc_fifo_0_out_endofpacket),                //          .endofpacket
		.data_out_data           (cpadderrouter_0_data_out_data),            //  data_out.data
		.data_out_valid          (cpadderrouter_0_data_out_valid),           //          .valid
		.data_out_error          (cpadderrouter_0_data_out_error),           //          .error
		.data_out_endofpacket    (cpadderrouter_0_data_out_endofpacket),     //          .endofpacket
		.data_out_startofpacket  (cpadderrouter_0_data_out_startofpacket)    //          .startofpacket
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (22),
		.FIFO_DEPTH          (32768),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (1),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sc_fifo_0 (
		.clk               (clk_clk),                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),           // clk_reset.reset
		.csr_address       (),                                         //       csr.address
		.csr_read          (),                                         //          .read
		.csr_write         (),                                         //          .write
		.csr_readdata      (),                                         //          .readdata
		.csr_writedata     (),                                         //          .writedata
		.in_data           (avalon_st_demux_0_aso_out1_data),          //        in.data
		.in_valid          (avalon_st_demux_0_aso_out1_valid),         //          .valid
		.in_ready          (avalon_st_demux_0_aso_out1_ready),         //          .ready
		.in_startofpacket  (avalon_st_demux_0_aso_out1_startofpacket), //          .startofpacket
		.in_endofpacket    (avalon_st_demux_0_aso_out1_endofpacket),   //          .endofpacket
		.out_data          (sc_fifo_0_out_data),                       //       out.data
		.out_valid         (sc_fifo_0_out_valid),                      //          .valid
		.out_ready         (sc_fifo_0_out_ready),                      //          .ready
		.out_startofpacket (sc_fifo_0_out_startofpacket),              //          .startofpacket
		.out_endofpacket   (sc_fifo_0_out_endofpacket),                //          .endofpacket
		.almost_full_data  (),                                         // (terminated)
		.almost_empty_data (),                                         // (terminated)
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.in_error          (1'b0),                                     // (terminated)
		.out_error         (),                                         // (terminated)
		.in_channel        (1'b0),                                     // (terminated)
		.out_channel       ()                                          // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
