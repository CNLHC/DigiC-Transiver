// DigiCQSysTop.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module DigiCQSysTop (
		input  wire        global_reset_reset_n,                    //              global_reset.reset_n
		output wire        pll_0_locked_export,                     //              pll_0_locked.export
		output wire        pll_0_outclk_1_clk,                      //            pll_0_outclk_1.clk
		output wire        pll_0_outclk_10_clk,                     //           pll_0_outclk_10.clk
		output wire        pll_0_outclk_120_clk,                    //          pll_0_outclk_120.clk
		output wire        pll_0_outclk_20_clk,                     //           pll_0_outclk_20.clk
		input  wire        pll_0_refclk_clk,                        //              pll_0_refclk.clk
		output wire [32:0] qam_modulation_0_aso_out0_data,          // qam_modulation_0_aso_out0.data
		input  wire        qam_modulation_0_aso_out0_ready,         //                          .ready
		output wire        qam_modulation_0_aso_out0_valid,         //                          .valid
		output wire        qam_modulation_0_aso_out0_empty,         //                          .empty
		output wire        qam_modulation_0_aso_out0_endofpacket,   //                          .endofpacket
		output wire        qam_modulation_0_aso_out0_startofpacket, //                          .startofpacket
		input  wire        qsys_clkin_clk,                          //                qsys_clkin.clk
		input  wire        spislave_0_export_0_mosi,                //       spislave_0_export_0.mosi
		input  wire        spislave_0_export_0_nss,                 //                          .nss
		inout  wire        spislave_0_export_0_miso,                //                          .miso
		input  wire        spislave_0_export_0_sclk                 //                          .sclk
	);

	DigiCQSysTop_DigiCQSys_0 digicqsys_0 (
		.global_reset_reset_n                    (global_reset_reset_n),                    //              global_reset.reset_n
		.pll_0_locked_export                     (pll_0_locked_export),                     //              pll_0_locked.export
		.pll_0_outclk_1_clk                      (pll_0_outclk_1_clk),                      //            pll_0_outclk_1.clk
		.pll_0_outclk_10_clk                     (pll_0_outclk_10_clk),                     //           pll_0_outclk_10.clk
		.pll_0_outclk_120_clk                    (pll_0_outclk_120_clk),                    //          pll_0_outclk_120.clk
		.pll_0_outclk_20_clk                     (pll_0_outclk_20_clk),                     //           pll_0_outclk_20.clk
		.pll_0_refclk_clk                        (pll_0_refclk_clk),                        //              pll_0_refclk.clk
		.qam_modulation_0_aso_out0_data          (qam_modulation_0_aso_out0_data),          // qam_modulation_0_aso_out0.data
		.qam_modulation_0_aso_out0_ready         (qam_modulation_0_aso_out0_ready),         //                          .ready
		.qam_modulation_0_aso_out0_valid         (qam_modulation_0_aso_out0_valid),         //                          .valid
		.qam_modulation_0_aso_out0_empty         (qam_modulation_0_aso_out0_empty),         //                          .empty
		.qam_modulation_0_aso_out0_endofpacket   (qam_modulation_0_aso_out0_endofpacket),   //                          .endofpacket
		.qam_modulation_0_aso_out0_startofpacket (qam_modulation_0_aso_out0_startofpacket), //                          .startofpacket
		.qsys_clkin_clk                          (qsys_clkin_clk),                          //                qsys_clkin.clk
		.spislave_0_export_0_mosi                (spislave_0_export_0_mosi),                //       spislave_0_export_0.mosi
		.spislave_0_export_0_nss                 (spislave_0_export_0_nss),                 //                          .nss
		.spislave_0_export_0_miso                (spislave_0_export_0_miso),                //                          .miso
		.spislave_0_export_0_sclk                (spislave_0_export_0_sclk)                 //                          .sclk
	);

endmodule
